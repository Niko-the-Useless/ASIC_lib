magic
tech scmos
timestamp 1742802875
<< checkpaint >>
rect 16 -27 34 -13
<< pwell >>
rect 17 -26 33 -16
<< polysilicon >>
rect 24 -18 26 -17
rect 24 -27 26 -24
<< ndiffusion >>
rect 17 -19 24 -18
rect 20 -23 24 -19
rect 17 -24 24 -23
rect 26 -19 33 -18
rect 26 -23 30 -19
rect 26 -24 33 -23
<< ntransistor >>
rect 24 -24 26 -18
<< polycontact >>
rect 23 -17 27 -13
<< ndcontact >>
rect 16 -23 20 -19
rect 30 -23 34 -19
<< labels >>
rlabel ndcontact 16 -23 20 -19 1 source
rlabel ndcontact 30 -23 34 -19 7 drain
rlabel polycontact 23 -17 27 -13 1 gate
<< end >>
