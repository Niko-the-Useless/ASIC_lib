magic
tech scmos
timestamp 1748381547
<< pwell >>
rect -140 -32 -70 -22
<< nwell >>
rect -140 -18 -70 -8
<< polysilicon >>
rect -135 -12 -133 -2
rect -127 -12 -125 -2
rect -119 -12 -117 -2
rect -111 -12 -109 -2
rect -103 -12 -101 -2
rect -95 -12 -93 -2
rect -87 -12 -85 -2
rect -79 -12 -77 -2
rect -135 -25 -133 -15
rect -127 -25 -125 -15
rect -119 -25 -117 -15
rect -111 -25 -109 -15
rect -103 -25 -101 -15
rect -95 -25 -93 -15
rect -87 -25 -85 -15
rect -79 -25 -77 -15
rect -135 -31 -133 -28
rect -127 -31 -125 -28
rect -119 -31 -117 -28
rect -111 -31 -109 -28
rect -103 -31 -101 -28
rect -95 -31 -93 -28
rect -87 -31 -85 -28
rect -79 -31 -77 -28
<< ndiffusion >>
rect -136 -28 -135 -25
rect -133 -28 -127 -25
rect -125 -28 -119 -25
rect -117 -28 -111 -25
rect -109 -28 -103 -25
rect -101 -28 -95 -25
rect -93 -28 -87 -25
rect -85 -28 -79 -25
rect -77 -28 -76 -25
rect -72 -28 -70 -25
<< pdiffusion >>
rect -136 -15 -135 -12
rect -133 -15 -132 -12
rect -128 -15 -127 -12
rect -125 -15 -124 -12
rect -120 -15 -119 -12
rect -117 -15 -116 -12
rect -112 -15 -111 -12
rect -109 -15 -108 -12
rect -104 -15 -103 -12
rect -101 -15 -100 -12
rect -96 -15 -95 -12
rect -93 -15 -92 -12
rect -88 -15 -87 -12
rect -85 -15 -84 -12
rect -80 -15 -79 -12
rect -77 -15 -76 -12
rect -72 -15 -70 -12
<< metal1 >>
rect -143 -8 -70 -5
rect -140 -11 -136 -8
rect -124 -11 -120 -8
rect -108 -11 -104 -8
rect -92 -11 -88 -8
rect -76 -11 -72 -8
rect -132 -18 -128 -15
rect -116 -18 -112 -15
rect -100 -18 -96 -15
rect -84 -18 -80 -15
rect -136 -22 -65 -18
rect -76 -25 -72 -22
rect -140 -32 -136 -29
rect -143 -35 -70 -32
<< ntransistor >>
rect -135 -28 -133 -25
rect -127 -28 -125 -25
rect -119 -28 -117 -25
rect -111 -28 -109 -25
rect -103 -28 -101 -25
rect -95 -28 -93 -25
rect -87 -28 -85 -25
rect -79 -28 -77 -25
<< ptransistor >>
rect -135 -15 -133 -12
rect -127 -15 -125 -12
rect -119 -15 -117 -12
rect -111 -15 -109 -12
rect -103 -15 -101 -12
rect -95 -15 -93 -12
rect -87 -15 -85 -12
rect -79 -15 -77 -12
<< polycontact >>
rect -136 -2 -132 2
rect -128 -2 -124 2
rect -120 -2 -116 2
rect -112 -2 -108 2
rect -104 -2 -100 2
rect -96 -2 -92 2
rect -88 -2 -84 2
rect -80 -2 -76 2
<< ndcontact >>
rect -140 -29 -136 -25
rect -76 -29 -72 -25
<< pdcontact >>
rect -140 -15 -136 -11
rect -132 -15 -128 -11
rect -124 -15 -120 -11
rect -116 -15 -112 -11
rect -108 -15 -104 -11
rect -100 -15 -96 -11
rect -92 -15 -88 -11
rect -84 -15 -80 -11
rect -76 -15 -72 -11
<< labels >>
rlabel metal1 -143 -35 -70 -32 1 Gnd
rlabel metal1 -143 -8 -70 -5 1 Vdd
rlabel polysilicon -135 -12 -133 -2 1 A
rlabel polysilicon -127 -12 -125 -2 1 B
rlabel metal1 -136 -22 -65 -18 1 Y
<< end >>
