magic
tech scmos
timestamp 1750012542
<< metal1 >>
rect -10 225 9 229
rect -40 199 -36 205
rect -40 195 -33 199
rect -25 177 -21 184
rect -25 166 -21 173
rect -40 155 -36 161
rect -40 151 -33 155
rect -10 124 -6 225
rect 19 210 44 214
rect -3 194 9 198
rect -3 177 1 194
rect 1 173 52 177
rect -3 156 1 173
rect -3 152 9 156
rect 19 136 44 140
rect -10 120 9 124
rect 66 -8 162 -4
rect 166 -8 290 -4
rect 294 -8 416 -4
rect 420 -8 542 -4
rect 546 -8 668 -4
rect 672 -8 681 -4
rect 66 -16 146 -12
rect 150 -16 252 -12
rect 256 -16 378 -12
rect 382 -16 504 -12
rect 508 -16 630 -12
rect 634 -16 681 -12
rect 66 -24 82 -20
rect 86 -24 227 -20
rect 231 -24 353 -20
rect 357 -24 479 -20
rect 483 -24 605 -20
rect 609 -24 681 -20
rect 70 -32 189 -28
rect 193 -32 315 -28
rect 319 -32 441 -28
rect 445 -32 567 -28
rect 571 -32 681 -28
rect 156 -47 176 -43
rect 8 -92 23 -88
rect 152 -92 166 -88
rect 162 -138 166 -92
rect 172 -111 176 -47
rect 172 -114 193 -111
rect 162 -142 191 -138
<< metal2 >>
rect 5 310 19 314
rect 5 252 9 310
rect 27 260 31 286
rect 27 256 48 260
rect 5 248 40 252
rect -33 210 2 214
rect -33 199 -29 210
rect -21 195 20 199
rect -21 173 -3 177
rect -21 151 20 155
rect -33 140 -29 151
rect -33 136 2 140
rect 36 -28 40 248
rect 44 214 48 256
rect 52 177 56 263
rect 4 -32 40 -28
rect 4 -88 8 -32
rect 44 -36 48 136
rect 26 -40 48 -36
rect 26 -71 30 -40
rect 52 -47 56 173
rect 66 -44 70 -32
rect 82 -44 86 -24
rect 146 -44 150 -16
rect 162 -44 166 -8
rect 181 -40 185 0
rect 189 -61 193 -32
rect 197 -40 201 8
rect 219 -40 223 16
rect 227 -61 231 -24
rect 235 -40 239 24
rect 244 -40 248 32
rect 252 -61 256 -16
rect 260 -40 264 40
rect 282 -40 286 48
rect 290 -61 294 -8
rect 298 -40 302 56
rect 317 24 321 64
rect 307 20 321 24
rect 307 -40 311 20
rect 335 16 339 72
rect 323 12 339 16
rect 315 -61 319 -32
rect 323 -40 327 12
rect 345 -40 349 80
rect 353 -61 357 -24
rect 361 -40 365 88
rect 370 -40 374 96
rect 378 -61 382 -16
rect 386 -40 390 104
rect 402 56 406 112
rect 402 52 412 56
rect 408 -40 412 52
rect 416 -61 420 -8
rect 424 -40 428 121
rect 433 -40 437 128
rect 441 -61 445 -32
rect 449 -40 453 136
rect 461 72 465 144
rect 482 80 486 152
rect 500 80 504 160
rect 482 76 491 80
rect 461 68 475 72
rect 471 -40 475 68
rect 479 -61 483 -24
rect 487 -40 491 76
rect 496 76 504 80
rect 496 -40 500 76
rect 504 -61 508 -16
rect 512 -40 516 168
rect 534 -40 538 176
rect 545 88 549 184
rect 564 88 568 192
rect 580 96 584 200
rect 545 84 554 88
rect 542 -61 546 -8
rect 550 -40 554 84
rect 559 84 568 88
rect 575 92 584 96
rect 559 -40 563 84
rect 567 -61 571 -32
rect 575 -40 579 92
rect 597 -40 601 208
rect 605 -61 609 -24
rect 613 -40 617 216
rect 622 -40 626 225
rect 644 104 648 232
rect 638 100 648 104
rect 630 -61 634 -16
rect 638 -40 642 100
rect 660 -40 664 240
rect 668 -61 672 -8
rect 676 -40 680 248
<< m2contact >>
rect 19 310 23 314
rect 52 263 56 267
rect 676 248 680 252
rect 660 240 664 244
rect 644 232 648 236
rect 622 225 626 229
rect -33 195 -29 199
rect -25 195 -21 199
rect -25 173 -21 177
rect -33 151 -29 155
rect -25 151 -21 155
rect 613 216 617 220
rect 2 210 6 214
rect 44 210 48 214
rect 597 208 601 212
rect 580 200 584 204
rect 564 192 568 196
rect 545 184 549 188
rect -3 173 1 177
rect 52 173 56 177
rect 534 176 538 180
rect 512 168 516 172
rect 500 160 504 164
rect 482 152 486 156
rect 461 144 465 148
rect 2 136 6 140
rect 44 136 48 140
rect 449 136 453 140
rect 433 128 437 132
rect 424 121 428 125
rect 402 112 406 116
rect 386 104 390 108
rect 370 96 374 100
rect 361 88 365 92
rect 345 80 349 84
rect 335 72 339 76
rect 317 64 321 68
rect 298 56 302 60
rect 282 48 286 52
rect 260 40 264 44
rect 244 32 248 36
rect 235 24 239 28
rect 219 16 223 20
rect 197 8 201 12
rect 181 0 185 4
rect 162 -8 166 -4
rect 290 -8 294 -4
rect 416 -8 420 -4
rect 542 -8 546 -4
rect 668 -8 672 -4
rect 146 -16 150 -12
rect 252 -16 256 -12
rect 378 -16 382 -12
rect 504 -16 508 -12
rect 630 -16 634 -12
rect 82 -24 86 -20
rect 227 -24 231 -20
rect 353 -24 357 -20
rect 479 -24 483 -20
rect 605 -24 609 -20
rect 66 -32 70 -28
rect 189 -32 193 -28
rect 315 -32 319 -28
rect 441 -32 445 -28
rect 567 -32 571 -28
rect 4 -92 8 -88
use inverter  inverter_0
timestamp 1749982892
transform 1 0 -10 0 1 200
box -22 -20 -9 14
use inverter  inverter_1
timestamp 1749982892
transform 1 0 -10 0 -1 150
box -22 -20 -9 14
use mux  mux_0
timestamp 1748844171
transform 1 0 5 0 1 212
box 0 -32 18 32
use mux  mux_1
timestamp 1748844171
transform 1 0 5 0 -1 138
box 0 -32 18 32
use nandArr  nandArr_0
timestamp 1749993027
transform 1 0 180 0 -1 -36
box 0 0 501 106
use shiftData2  shiftData2_0
timestamp 1749984423
transform 1 0 -1 0 -1 -36
box 0 0 1 1
use shiftData32  shiftData32_0
timestamp 1749990304
transform 1 0 -1308 0 1 -128
box 1308 128 2625 444
use shiftreg2  shiftreg2_0
timestamp 1749982892
transform 1 0 -1 0 -1 -43
box 0 -7 167 53
<< labels >>
rlabel metal1 -40 195 -36 205 3 progEN
rlabel metal1 -40 151 -36 161 3 dataEN
<< end >>
