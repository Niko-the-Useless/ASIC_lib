magic
tech scmos
timestamp 1749993027
<< pwell >>
rect -7 -58 29 -48
<< nwell >>
rect -7 -44 29 -34
<< polysilicon >>
rect -2 -38 0 -20
rect 6 -38 8 -20
rect 14 -38 16 -20
rect 22 -38 24 -20
rect -2 -51 0 -41
rect 6 -51 8 -41
rect 14 -51 16 -41
rect 22 -51 24 -41
rect -2 -57 0 -54
rect 6 -57 8 -54
rect 14 -57 16 -54
rect 22 -57 24 -54
<< ndiffusion >>
rect -3 -54 -2 -51
rect 0 -54 6 -51
rect 8 -54 14 -51
rect 16 -54 22 -51
rect 24 -54 25 -51
<< pdiffusion >>
rect -3 -41 -2 -38
rect 0 -41 1 -38
rect 5 -41 6 -38
rect 8 -41 9 -38
rect 13 -41 14 -38
rect 16 -41 17 -38
rect 21 -41 22 -38
rect 24 -41 25 -38
<< metal1 >>
rect 25 -28 43 -24
rect 25 -30 29 -28
rect -7 -34 29 -30
rect 39 -33 43 -28
rect -7 -37 -3 -34
rect 9 -37 13 -34
rect 25 -37 29 -34
rect 1 -44 5 -41
rect 17 -44 21 -41
rect -7 -48 29 -44
rect 25 -51 29 -48
rect -7 -58 -3 -55
rect -7 -62 29 -58
<< ntransistor >>
rect -2 -54 0 -51
rect 6 -54 8 -51
rect 14 -54 16 -51
rect 22 -54 24 -51
<< ptransistor >>
rect -2 -41 0 -38
rect 6 -41 8 -38
rect 14 -41 16 -38
rect 22 -41 24 -38
<< polycontact >>
rect -3 -20 1 -16
rect 5 -20 9 -16
rect 13 -20 17 -16
rect 21 -20 25 -16
<< ndcontact >>
rect -7 -55 -3 -51
rect 25 -55 29 -51
<< pdcontact >>
rect -7 -41 -3 -37
rect 1 -41 5 -37
rect 9 -41 13 -37
rect 17 -41 21 -37
rect 25 -41 29 -37
<< labels >>
rlabel metal1 -7 -48 29 -44 1 Y
<< end >>
