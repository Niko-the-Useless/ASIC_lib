magic
tech scmos
timestamp 1745822104
<< pwell >>
rect -1 10 9 26
rect 50 5 60 21
rect -1 -16 9 0
rect -1 -93 9 -77
rect 50 -98 60 -82
rect -1 -119 9 -103
<< nwell >>
rect -1 44 9 62
rect 22 44 32 62
rect 50 37 60 55
rect -1 -59 9 -41
rect 22 -59 32 -41
rect 50 -66 60 -48
<< polysilicon >>
rect 0 52 1 54
rect 7 52 10 54
rect 23 52 24 54
rect 30 52 33 54
rect 51 45 52 47
rect 58 45 61 47
rect 0 17 1 19
rect 7 17 10 19
rect 51 12 52 14
rect 58 12 61 14
rect 0 -9 1 -7
rect 7 -9 10 -7
rect 0 -51 1 -49
rect 7 -51 10 -49
rect 23 -51 24 -49
rect 30 -51 33 -49
rect 51 -58 52 -56
rect 58 -58 61 -56
rect 0 -86 1 -84
rect 7 -86 10 -84
rect 51 -91 52 -89
rect 58 -91 61 -89
rect 0 -112 1 -110
rect 7 -112 10 -110
<< ndiffusion >>
rect 1 23 2 26
rect 6 23 7 26
rect 1 19 7 23
rect 52 18 53 21
rect 57 18 58 21
rect 1 13 7 17
rect 1 10 2 13
rect 6 10 7 13
rect 52 14 58 18
rect 52 8 58 12
rect 52 5 53 8
rect 57 5 58 8
rect 1 -3 2 0
rect 6 -3 7 0
rect 1 -7 7 -3
rect 1 -13 7 -9
rect 1 -16 2 -13
rect 6 -16 7 -13
rect 1 -80 2 -77
rect 6 -80 7 -77
rect 1 -84 7 -80
rect 52 -85 53 -82
rect 57 -85 58 -82
rect 1 -90 7 -86
rect 1 -93 2 -90
rect 6 -93 7 -90
rect 52 -89 58 -85
rect 52 -95 58 -91
rect 52 -98 53 -95
rect 57 -98 58 -95
rect 1 -106 2 -103
rect 6 -106 7 -103
rect 1 -110 7 -106
rect 1 -116 7 -112
rect 1 -119 2 -116
rect 6 -119 7 -116
<< pdiffusion >>
rect 1 58 2 61
rect 6 58 7 61
rect 1 54 7 58
rect 24 58 25 61
rect 29 58 30 61
rect 1 48 7 52
rect 24 54 30 58
rect 1 45 2 48
rect 6 45 7 48
rect 24 48 30 52
rect 52 51 53 54
rect 57 51 58 54
rect 24 45 25 48
rect 29 45 30 48
rect 52 47 58 51
rect 52 41 58 45
rect 52 38 53 41
rect 57 38 58 41
rect 1 -45 2 -42
rect 6 -45 7 -42
rect 1 -49 7 -45
rect 24 -45 25 -42
rect 29 -45 30 -42
rect 1 -55 7 -51
rect 24 -49 30 -45
rect 1 -58 2 -55
rect 6 -58 7 -55
rect 24 -55 30 -51
rect 52 -52 53 -49
rect 57 -52 58 -49
rect 24 -58 25 -55
rect 29 -58 30 -55
rect 52 -56 58 -52
rect 52 -62 58 -58
rect 52 -65 53 -62
rect 57 -65 58 -62
<< metal1 >>
rect 53 69 104 73
rect -22 65 57 69
rect 2 62 6 65
rect 25 62 29 65
rect 53 55 57 65
rect -10 51 -4 55
rect 14 51 19 55
rect -10 41 -6 51
rect -22 37 -6 41
rect -10 20 -6 37
rect 2 41 6 44
rect 25 41 29 44
rect 41 44 47 48
rect 41 41 45 44
rect 81 41 106 45
rect 2 37 45 41
rect 2 27 6 37
rect -10 16 -4 20
rect 41 15 45 37
rect 53 31 57 37
rect 81 31 85 41
rect 53 27 85 31
rect 53 22 57 27
rect 41 11 47 15
rect 2 1 6 9
rect -9 -10 -4 -6
rect 2 -19 6 -17
rect 53 -15 57 4
rect 53 -19 100 -15
rect -22 -23 57 -19
rect -22 -38 57 -34
rect 2 -41 6 -38
rect 25 -41 29 -38
rect 53 -42 100 -38
rect 53 -48 57 -42
rect -10 -52 -4 -48
rect 14 -52 19 -48
rect -10 -62 -6 -52
rect -22 -66 -6 -62
rect -10 -83 -6 -66
rect 2 -62 6 -59
rect 25 -62 29 -59
rect 41 -59 47 -55
rect 41 -62 45 -59
rect 2 -66 45 -62
rect 2 -76 6 -66
rect -10 -87 -4 -83
rect 41 -88 45 -66
rect 53 -72 57 -66
rect 53 -76 82 -72
rect 53 -81 57 -76
rect 78 -87 82 -76
rect 41 -92 47 -88
rect 2 -102 6 -94
rect -9 -113 -4 -109
rect 2 -122 6 -120
rect 53 -122 57 -99
rect -22 -126 57 -122
rect 53 -130 104 -126
<< metal2 >>
rect -14 51 13 55
rect -14 20 -10 51
rect -22 16 -10 20
rect -14 -10 -10 16
rect -14 -52 13 -48
rect -14 -83 -10 -52
rect -22 -87 -10 -83
rect -14 -113 -10 -87
rect 82 -91 104 -87
<< ntransistor >>
rect 1 17 7 19
rect 52 12 58 14
rect 1 -9 7 -7
rect 1 -86 7 -84
rect 52 -91 58 -89
rect 1 -112 7 -110
<< ptransistor >>
rect 1 52 7 54
rect 24 52 30 54
rect 52 45 58 47
rect 1 -51 7 -49
rect 24 -51 30 -49
rect 52 -58 58 -56
<< polycontact >>
rect -4 51 0 55
rect 19 51 23 55
rect 47 44 51 48
rect -4 16 0 20
rect 47 11 51 15
rect -4 -10 0 -6
rect -4 -52 0 -48
rect 19 -52 23 -48
rect 47 -59 51 -55
rect -4 -87 0 -83
rect 47 -92 51 -88
rect -4 -113 0 -109
<< ndcontact >>
rect 2 23 6 27
rect 53 18 57 22
rect 2 9 6 13
rect 53 4 57 8
rect 2 -3 6 1
rect 2 -17 6 -13
rect 2 -80 6 -76
rect 53 -85 57 -81
rect 2 -94 6 -90
rect 53 -99 57 -95
rect 2 -106 6 -102
rect 2 -120 6 -116
<< pdcontact >>
rect 2 58 6 62
rect 25 58 29 62
rect 2 44 6 48
rect 53 51 57 55
rect 25 44 29 48
rect 53 37 57 41
rect 2 -45 6 -41
rect 25 -45 29 -41
rect 2 -59 6 -55
rect 53 -52 57 -48
rect 25 -59 29 -55
rect 53 -66 57 -62
<< m2contact >>
rect 78 -91 82 -87
<< pad >>
rect 13 51 19 55
rect -10 -10 -4 -6
rect 13 -52 19 -48
rect -10 -113 -4 -109
<< labels >>
rlabel metal1 -22 -126 -13 -122 3 Gnd
rlabel metal1 -22 -38 -13 -34 3 Vdd
rlabel metal1 -22 -23 -13 -19 3 Gnd
rlabel metal1 -22 65 -13 69 3 Vdd
rlabel metal1 -22 -66 -17 -62 3 CLK
rlabel metal2 -22 -87 -17 -83 3 RESET
rlabel metal2 -22 16 -17 20 3 CLK
rlabel metal1 -22 37 -17 41 3 SET
<< end >>
