magic
tech scmos
timestamp 1749937379
<< pwell >>
rect -140 -32 -120 -22
<< nwell >>
rect -140 -18 -120 -8
<< polysilicon >>
rect -135 -12 -133 -9
rect -127 -12 -125 -9
rect -135 -25 -133 -15
rect -127 -25 -125 -15
rect -135 -38 -133 -28
rect -127 -38 -125 -28
<< ndiffusion >>
rect -136 -28 -135 -25
rect -133 -28 -127 -25
rect -125 -28 -124 -25
<< pdiffusion >>
rect -136 -15 -135 -12
rect -133 -15 -132 -12
rect -128 -15 -127 -12
rect -125 -15 -124 -12
<< ntransistor >>
rect -135 -28 -133 -25
rect -127 -28 -125 -25
<< ptransistor >>
rect -135 -15 -133 -12
rect -127 -15 -125 -12
<< polycontact >>
rect -136 -42 -132 -38
rect -128 -42 -124 -38
<< ndcontact >>
rect -140 -29 -136 -25
rect -124 -29 -120 -25
<< pdcontact >>
rect -140 -15 -136 -11
rect -132 -15 -128 -11
rect -124 -15 -120 -11
<< end >>
