magic
tech scmos
timestamp 1748847516
<< pwell >>
rect 2 -30 13 -11
<< nwell >>
rect 2 -1 13 18
<< polysilicon >>
rect 4 11 7 13
rect 11 11 13 13
rect 4 4 7 6
rect 11 4 13 6
rect 4 -18 7 -16
rect 11 -18 13 -16
rect 4 -25 7 -23
rect 11 -25 13 -23
<< ndiffusion >>
rect 7 -16 11 -15
rect 7 -23 11 -18
rect 7 -26 11 -25
<< pdiffusion >>
rect 7 13 11 14
rect 7 6 11 11
rect 7 3 11 4
<< metal1 >>
rect -11 10 0 14
rect -11 -22 -8 10
rect -1 3 0 7
rect 7 -11 11 -1
rect -1 -19 0 -15
rect -11 -26 0 -22
<< ntransistor >>
rect 7 -18 11 -16
rect 7 -25 11 -23
<< ptransistor >>
rect 7 11 11 13
rect 7 4 11 6
<< polycontact >>
rect 0 10 4 14
rect 0 3 4 7
rect 0 -19 4 -15
rect 0 -26 4 -22
<< ndcontact >>
rect 7 -15 11 -11
rect 7 -30 11 -26
<< pdcontact >>
rect 7 14 11 18
rect 7 -1 11 3
<< m2contact >>
rect -5 3 -1 7
rect -5 -19 -1 -15
<< end >>
