magic
tech scmos
timestamp 1747033067
<< pwell >>
rect 99 -91 115 -81
rect 133 -91 149 -81
rect -150 -118 -134 -108
rect -150 -148 -134 -138
rect 27 -145 37 -129
rect 53 -145 63 -129
rect 42 -174 52 -158
<< nwell >>
rect -150 -96 -134 -86
rect 27 -113 37 -97
rect 53 -113 63 -97
rect 99 -107 115 -97
rect 133 -107 149 -97
rect -150 -170 -134 -160
<< polysilicon >>
rect 106 -83 108 -82
rect 140 -83 142 -82
rect -143 -88 -141 -87
rect 106 -91 108 -89
rect 140 -91 142 -89
rect -143 -110 -141 -94
rect -143 -119 -141 -116
rect -129 -124 -125 -100
rect 106 -99 108 -97
rect 140 -99 142 -97
rect 26 -106 29 -104
rect 35 -106 36 -104
rect 54 -106 55 -104
rect 61 -106 64 -104
rect 106 -106 108 -105
rect 140 -106 142 -105
rect -157 -132 -125 -124
rect -143 -140 -141 -137
rect -143 -162 -141 -146
rect -129 -156 -125 -132
rect 82 -135 86 -118
rect 28 -138 29 -136
rect 35 -138 38 -136
rect 52 -138 55 -136
rect 61 -138 62 -136
rect 78 -139 86 -135
rect 82 -156 86 -139
rect 43 -167 44 -165
rect 50 -167 53 -165
rect -143 -169 -141 -168
<< ndiffusion >>
rect 99 -84 106 -83
rect 102 -88 106 -84
rect 99 -89 106 -88
rect 108 -84 115 -83
rect 133 -84 140 -83
rect 108 -88 112 -84
rect 136 -88 140 -84
rect 108 -89 115 -88
rect 133 -89 140 -88
rect 142 -84 149 -83
rect 142 -88 146 -84
rect 142 -89 149 -88
rect -150 -111 -143 -110
rect -147 -115 -143 -111
rect -150 -116 -143 -115
rect -141 -111 -134 -110
rect -141 -115 -137 -111
rect -141 -116 -134 -115
rect -150 -141 -143 -140
rect -147 -145 -143 -141
rect -150 -146 -143 -145
rect -141 -141 -134 -140
rect -141 -145 -137 -141
rect -141 -146 -134 -145
rect 29 -132 30 -129
rect 34 -132 35 -129
rect 29 -136 35 -132
rect 55 -132 56 -129
rect 60 -132 61 -129
rect 55 -136 61 -132
rect 29 -142 35 -138
rect 29 -145 30 -142
rect 34 -145 35 -142
rect 55 -142 61 -138
rect 55 -145 56 -142
rect 60 -145 61 -142
rect 44 -161 45 -158
rect 49 -161 50 -158
rect 44 -165 50 -161
rect 44 -171 50 -167
rect 44 -174 45 -171
rect 49 -174 50 -171
<< pdiffusion >>
rect -150 -89 -143 -88
rect -147 -93 -143 -89
rect -150 -94 -143 -93
rect -141 -89 -134 -88
rect -141 -93 -137 -89
rect -141 -94 -134 -93
rect 29 -100 30 -97
rect 34 -100 35 -97
rect 29 -104 35 -100
rect 55 -100 56 -97
rect 60 -100 61 -97
rect 99 -100 106 -99
rect 29 -110 35 -106
rect 55 -104 61 -100
rect 102 -104 106 -100
rect 99 -105 106 -104
rect 108 -100 115 -99
rect 133 -100 140 -99
rect 108 -104 112 -100
rect 136 -104 140 -100
rect 108 -105 115 -104
rect 133 -105 140 -104
rect 142 -100 149 -99
rect 142 -104 146 -100
rect 142 -105 149 -104
rect 29 -113 30 -110
rect 34 -113 35 -110
rect 55 -110 61 -106
rect 55 -113 56 -110
rect 60 -113 61 -110
rect -150 -163 -143 -162
rect -147 -167 -143 -163
rect -150 -168 -143 -167
rect -141 -163 -134 -162
rect -141 -167 -137 -163
rect -141 -168 -134 -167
<< metal1 >>
rect 43 -87 47 -81
rect -137 -111 -133 -93
rect 30 -91 60 -87
rect 30 -96 34 -91
rect 56 -96 60 -91
rect 98 -92 102 -88
rect 82 -96 102 -92
rect 40 -107 50 -103
rect 30 -118 34 -114
rect 43 -118 47 -107
rect 30 -122 47 -118
rect 82 -114 86 -96
rect 98 -100 102 -96
rect 112 -92 116 -88
rect 132 -92 136 -88
rect 112 -96 136 -92
rect 112 -100 116 -96
rect 119 -113 124 -96
rect 132 -100 136 -96
rect 146 -92 150 -88
rect 146 -96 163 -92
rect 146 -100 150 -96
rect 153 -113 158 -96
rect 56 -118 82 -114
rect 30 -128 34 -122
rect 56 -128 60 -118
rect 16 -139 24 -135
rect 66 -139 74 -135
rect -137 -163 -133 -145
rect 34 -146 56 -142
rect 45 -157 49 -146
rect 55 -160 82 -156
rect 97 -159 126 -113
rect 131 -159 160 -113
rect 29 -168 39 -164
rect 29 -179 33 -168
rect 45 -179 49 -175
rect 55 -179 59 -160
rect 82 -162 86 -160
rect 82 -166 109 -162
rect 113 -166 143 -162
rect 16 -183 59 -179
<< metal2 >>
rect 105 -110 109 -74
rect 139 -110 143 -74
rect 97 -162 126 -116
rect 97 -164 109 -162
rect 113 -164 126 -162
rect 131 -162 160 -116
rect 131 -164 143 -162
rect 147 -164 160 -162
<< ntransistor >>
rect 106 -89 108 -83
rect 140 -89 142 -83
rect -143 -116 -141 -110
rect -143 -146 -141 -140
rect 29 -138 35 -136
rect 55 -138 61 -136
rect 44 -167 50 -165
<< ptransistor >>
rect -143 -94 -141 -88
rect 29 -106 35 -104
rect 55 -106 61 -104
rect 106 -105 108 -99
rect 140 -105 142 -99
rect -143 -168 -141 -162
<< polycontact >>
rect 105 -82 109 -78
rect 139 -82 143 -78
rect -144 -87 -140 -83
rect -133 -104 -129 -100
rect 36 -107 40 -103
rect 50 -107 54 -103
rect 105 -110 109 -106
rect 139 -110 143 -106
rect 82 -118 86 -114
rect -133 -156 -129 -152
rect 24 -139 28 -135
rect 62 -139 66 -135
rect 74 -139 78 -135
rect 82 -160 86 -156
rect 39 -168 43 -164
rect -144 -173 -140 -169
<< ndcontact >>
rect 98 -88 102 -84
rect 112 -88 116 -84
rect 132 -88 136 -84
rect 146 -88 150 -84
rect -151 -115 -147 -111
rect -137 -115 -133 -111
rect -151 -145 -147 -141
rect -137 -145 -133 -141
rect 30 -132 34 -128
rect 56 -132 60 -128
rect 30 -146 34 -142
rect 56 -146 60 -142
rect 45 -161 49 -157
rect 45 -175 49 -171
<< pdcontact >>
rect -151 -93 -147 -89
rect -137 -93 -133 -89
rect 30 -100 34 -96
rect 56 -100 60 -96
rect 98 -104 102 -100
rect 112 -104 116 -100
rect 132 -104 136 -100
rect 146 -104 150 -100
rect 30 -114 34 -110
rect 56 -114 60 -110
rect -151 -167 -147 -163
rect -137 -167 -133 -163
<< m2contact >>
rect 109 -166 113 -162
rect 143 -166 147 -162
<< labels >>
rlabel metal1 16 -139 20 -135 3 In2
rlabel metal1 43 -85 47 -81 5 Vdd
rlabel metal1 16 -183 20 -179 2 Gnd
rlabel pdcontact -151 -93 -147 -89 3 vdd
rlabel polycontact -144 -87 -140 -83 1 in
rlabel pdcontact -151 -167 -147 -163 3 vdd
rlabel polycontact -144 -173 -140 -169 5 in
<< end >>
