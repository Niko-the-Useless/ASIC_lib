magic
tech scmos
timestamp 1748365915
<< metal1 >>
rect 12 75 16 82
rect 37 75 41 82
rect -1 64 72 68
rect -1 51 3 64
rect 29 56 53 60
rect 29 52 33 56
rect 49 52 53 56
rect 68 51 72 64
rect -12 37 -1 41
rect 3 37 12 41
rect 16 37 26 41
rect 29 37 37 41
rect 41 37 42 41
rect 49 37 68 41
rect 72 37 85 41
rect -1 22 3 27
rect -15 18 3 22
rect 12 7 16 37
rect 29 22 33 26
rect 49 22 53 26
rect 29 18 53 22
rect 68 18 72 27
rect 81 7 85 37
rect 12 3 85 7
<< metal2 >>
rect 12 41 16 71
rect 37 41 41 71
rect 3 14 68 18
<< m2contact >>
rect 12 71 16 75
rect 37 71 41 75
rect 12 37 16 41
rect 37 37 41 41
rect -1 14 3 18
rect 68 14 72 18
use inverter  inverter_0
timestamp 1748362390
transform 1 0 44 0 1 42
box -22 -20 -9 14
use inverter  inverter_1
timestamp 1748362390
transform 1 0 64 0 1 42
box -22 -20 -9 14
use transgate  transgate_0
timestamp 1748362827
transform 1 0 0 0 1 62
box -5 -39 7 -7
use transgate  transgate_1
timestamp 1748362827
transform 1 0 69 0 -1 16
box -5 -39 7 -7
<< labels >>
rlabel metal1 -12 37 -1 41 1 D
rlabel metal1 -15 18 3 22 1 NC
rlabel metal1 -1 64 72 68 5 CC
rlabel metal1 29 56 53 60 1 Vdd
rlabel metal1 29 18 53 22 1 Gnd
rlabel metal1 12 75 16 82 5 Q
rlabel metal1 37 75 41 82 5 NQ
<< end >>
