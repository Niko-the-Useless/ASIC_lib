magic
tech scmos
timestamp 1746427415
<< pwell >>
rect 5 -16 15 0
rect 31 -16 41 0
rect 20 -45 30 -29
<< nwell >>
rect 5 16 15 32
rect 31 16 41 32
<< polysilicon >>
rect 4 23 7 25
rect 13 23 14 25
rect 32 23 33 25
rect 39 23 42 25
rect 60 0 64 11
rect 60 -4 107 0
rect 6 -9 7 -7
rect 13 -9 16 -7
rect 30 -9 33 -7
rect 39 -9 40 -7
rect 56 -10 87 -6
rect 83 -12 87 -10
rect 103 -12 107 -4
rect 60 -16 107 -12
rect 60 -18 64 -16
rect 60 -22 107 -18
rect 103 -24 107 -22
rect 60 -27 107 -24
rect 64 -28 107 -27
rect 21 -38 22 -36
rect 28 -38 31 -36
<< ndiffusion >>
rect 7 -3 8 0
rect 12 -3 13 0
rect 7 -7 13 -3
rect 33 -3 34 0
rect 38 -3 39 0
rect 33 -7 39 -3
rect 7 -13 13 -9
rect 7 -16 8 -13
rect 12 -16 13 -13
rect 33 -13 39 -9
rect 33 -16 34 -13
rect 38 -16 39 -13
rect 22 -32 23 -29
rect 27 -32 28 -29
rect 22 -36 28 -32
rect 22 -42 28 -38
rect 22 -45 23 -42
rect 27 -45 28 -42
<< pdiffusion >>
rect 7 29 8 32
rect 12 29 13 32
rect 7 25 13 29
rect 33 29 34 32
rect 38 29 39 32
rect 7 19 13 23
rect 33 25 39 29
rect 7 16 8 19
rect 12 16 13 19
rect 33 19 39 23
rect 33 16 34 19
rect 38 16 39 19
<< metal1 >>
rect 21 42 25 48
rect 8 38 38 42
rect 8 33 12 38
rect 34 33 38 38
rect 18 22 28 26
rect 8 11 12 15
rect 21 11 25 22
rect 8 7 25 11
rect 34 11 60 15
rect 64 11 70 15
rect 8 1 12 7
rect 34 1 38 11
rect -6 -10 2 -6
rect 44 -10 52 -6
rect 12 -17 34 -13
rect 23 -28 27 -17
rect 7 -39 17 -35
rect 7 -50 11 -39
rect 23 -50 27 -46
rect 60 -50 64 -31
rect -6 -54 64 -50
<< ntransistor >>
rect 7 -9 13 -7
rect 33 -9 39 -7
rect 22 -38 28 -36
<< ptransistor >>
rect 7 23 13 25
rect 33 23 39 25
<< polycontact >>
rect 14 22 18 26
rect 28 22 32 26
rect 60 11 64 15
rect 2 -10 6 -6
rect 40 -10 44 -6
rect 52 -10 56 -6
rect 60 -31 64 -27
rect 17 -39 21 -35
<< ndcontact >>
rect 8 -3 12 1
rect 34 -3 38 1
rect 8 -17 12 -13
rect 34 -17 38 -13
rect 23 -32 27 -28
rect 23 -46 27 -42
<< pdcontact >>
rect 8 29 12 33
rect 34 29 38 33
rect 8 15 12 19
rect 34 15 38 19
<< labels >>
rlabel metal1 -6 -54 -2 -50 2 Gnd
rlabel metal1 -6 -10 -2 -6 3 In2
rlabel metal1 21 44 25 48 5 Vdd
rlabel metal1 70 11 74 15 7 Out
<< end >>
