magic
tech scmos
timestamp 1750012542
<< metal1 >>
rect -1 450 28 454
rect -1 446 3 450
rect -3 428 6 432
rect -3 423 1 428
rect 0 405 29 409
rect 0 401 4 405
rect -4 76 0 83
rect -4 72 5 76
rect 733 39 762 43
rect 680 35 692 39
rect 680 31 683 35
rect 733 32 737 39
rect 669 28 683 31
rect 822 19 826 25
rect 818 15 826 19
rect 670 0 687 4
rect 733 -2 737 6
rect 291 -8 695 -4
rect 699 -12 703 -4
rect 287 -16 413 -12
rect 417 -16 703 -12
rect 707 -20 711 -4
rect 287 -24 539 -20
rect 543 -24 711 -20
rect 715 -29 719 -4
rect 733 -6 764 -2
rect 287 -33 665 -29
rect 669 -33 719 -29
<< metal2 >>
rect 771 47 775 458
rect 762 43 775 47
rect 762 25 766 43
rect 287 -4 291 14
rect 413 -12 417 14
rect 539 -20 543 14
rect 665 -29 669 14
<< m2contact >>
rect 29 454 33 458
rect 287 14 291 18
rect 413 14 417 18
rect 539 14 543 18
rect 665 14 669 18
rect 287 -8 291 -4
rect 413 -16 417 -12
rect 539 -24 543 -20
rect 665 -33 669 -29
use and4  and4_0
timestamp 1749993027
transform 1 0 706 0 -1 -8
box -25 -47 33 0
use pla1stage  pla1stage_0
timestamp 1750012542
transform 1 0 2 0 1 142
box -40 -142 1317 316
use TSPCff  TSPCff_0
timestamp 1749982892
transform 1 0 767 0 -1 8
box -32 -35 55 14
<< labels >>
rlabel metal1 822 15 826 25 1 Y
rlabel metal1 -4 72 0 83 3 IN
rlabel metal1 -3 423 1 432 3 PROGRAM
rlabel metal1 -1 446 3 454 3 Vdd
rlabel metal1 0 401 4 409 1 Gnd
<< end >>
