magic
tech scmos
timestamp 1748253556
<< pwell >>
rect -139 -31 -101 -21
<< nwell >>
rect -139 -17 -101 -7
<< polysilicon >>
rect -134 -11 -132 -2
rect -126 -11 -124 -2
rect -118 -11 -116 -2
rect -110 -11 -108 -2
rect -134 -24 -132 -14
rect -126 -24 -124 -14
rect -118 -24 -116 -14
rect -110 -24 -108 -14
rect -134 -30 -132 -27
rect -126 -30 -124 -27
rect -118 -30 -116 -27
rect -110 -30 -108 -27
<< ndiffusion >>
rect -135 -27 -134 -24
rect -132 -27 -126 -24
rect -124 -27 -118 -24
rect -116 -27 -110 -24
rect -108 -27 -107 -24
rect -103 -27 -101 -24
<< pdiffusion >>
rect -135 -14 -134 -11
rect -132 -14 -131 -11
rect -127 -14 -126 -11
rect -124 -14 -123 -11
rect -119 -14 -118 -11
rect -116 -14 -115 -11
rect -111 -14 -110 -11
rect -108 -14 -107 -11
rect -103 -14 -101 -11
<< metal1 >>
rect -142 -7 -101 -4
rect -139 -10 -135 -7
rect -123 -10 -119 -7
rect -107 -10 -103 -7
rect -139 -31 -135 -28
rect -142 -34 -101 -31
<< metal2 >>
rect -131 -17 -127 -10
rect -115 -17 -111 -10
rect -139 -21 -97 -17
rect -107 -28 -103 -21
<< ntransistor >>
rect -134 -27 -132 -24
rect -126 -27 -124 -24
rect -118 -27 -116 -24
rect -110 -27 -108 -24
<< ptransistor >>
rect -134 -14 -132 -11
rect -126 -14 -124 -11
rect -118 -14 -116 -11
rect -110 -14 -108 -11
<< ndcontact >>
rect -139 -28 -135 -24
rect -107 -28 -103 -24
<< pdcontact >>
rect -139 -14 -135 -10
rect -131 -14 -127 -10
rect -123 -14 -119 -10
rect -115 -14 -111 -10
rect -107 -14 -103 -10
<< labels >>
rlabel metal1 -142 -7 -101 -4 5 Vdd
rlabel metal1 -142 -34 -101 -31 1 Gnd
rlabel polysilicon -134 -11 -132 -2 5 A
rlabel polysilicon -126 -11 -124 -2 5 B
rlabel polysilicon -118 -11 -116 -2 5 C
rlabel polysilicon -110 -11 -108 -2 5 D
rlabel metal2 -139 -21 -97 -17 1 Y
<< end >>
