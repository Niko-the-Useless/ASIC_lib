magic
tech scmos
timestamp 1749990304
<< metal1 >>
rect 1374 376 2625 380
rect 1374 368 2598 372
rect 2602 368 2625 372
rect 1374 360 2534 364
rect 2538 360 2625 364
rect 1374 352 2518 356
rect 2522 352 2625 356
rect 1374 344 2452 348
rect 2456 344 2625 348
rect 1374 336 2436 340
rect 2440 336 2625 340
rect 1374 328 2372 332
rect 2376 328 2625 332
rect 1374 320 2356 324
rect 2360 320 2625 324
rect 1374 312 2287 316
rect 2291 312 2625 316
rect 1374 304 2271 308
rect 2275 304 2625 308
rect 1374 296 2207 300
rect 2211 296 2625 300
rect 1374 288 2191 292
rect 2195 288 2625 292
rect 1374 280 2125 284
rect 2129 280 2625 284
rect 1374 272 2109 276
rect 2113 272 2625 276
rect 1374 264 2045 268
rect 2049 264 2625 268
rect 1374 256 2029 260
rect 2033 256 2625 260
rect 1374 248 1960 252
rect 1964 248 2625 252
rect 1374 240 1944 244
rect 1948 240 2625 244
rect 1374 232 1880 236
rect 1884 232 2625 236
rect 1374 224 1864 228
rect 1868 224 2625 228
rect 1374 216 1798 220
rect 1802 216 2625 220
rect 1374 208 1782 212
rect 1786 208 2625 212
rect 1374 200 1718 204
rect 1722 200 2625 204
rect 1374 192 1702 196
rect 1706 192 2625 196
rect 1374 184 1633 188
rect 1637 184 2625 188
rect 1374 176 1617 180
rect 1621 176 2625 180
rect 1374 168 1553 172
rect 1557 168 2625 172
rect 1374 160 1537 164
rect 1541 160 2625 164
rect 1374 152 1471 156
rect 1475 152 2625 156
rect 1374 144 1455 148
rect 1459 144 2625 148
rect 1374 136 1391 140
rect 1395 136 2625 140
rect 1374 128 1375 132
rect 1379 128 2625 132
<< metal2 >>
rect 1375 132 1379 388
rect 1391 140 1395 388
rect 1455 148 1459 388
rect 1471 156 1475 388
rect 1537 164 1541 388
rect 1553 172 1557 388
rect 1617 180 1621 388
rect 1633 188 1637 388
rect 1702 196 1706 388
rect 1718 204 1722 388
rect 1782 212 1786 388
rect 1798 220 1802 388
rect 1864 228 1868 388
rect 1880 236 1884 388
rect 1944 244 1948 388
rect 1960 252 1964 388
rect 2029 260 2033 388
rect 2045 268 2049 388
rect 2109 276 2113 399
rect 2125 284 2129 399
rect 2191 292 2195 419
rect 2207 300 2211 419
rect 2271 308 2275 392
rect 2287 316 2291 392
rect 2356 324 2360 392
rect 2372 332 2376 392
rect 2436 340 2440 392
rect 2452 348 2456 392
rect 2518 356 2522 392
rect 2534 364 2538 392
rect 2598 372 2602 392
rect 2614 376 2618 393
<< m2contact >>
rect 2598 368 2602 372
rect 2534 360 2538 364
rect 2518 352 2522 356
rect 2452 344 2456 348
rect 2436 336 2440 340
rect 2372 328 2376 332
rect 2356 320 2360 324
rect 2287 312 2291 316
rect 2271 304 2275 308
rect 2207 296 2211 300
rect 2191 288 2195 292
rect 2125 280 2129 284
rect 2109 272 2113 276
rect 2045 264 2049 268
rect 2029 256 2033 260
rect 1960 248 1964 252
rect 1944 240 1948 244
rect 1880 232 1884 236
rect 1864 224 1868 228
rect 1798 216 1802 220
rect 1782 208 1786 212
rect 1718 200 1722 204
rect 1702 192 1706 196
rect 1633 184 1637 188
rect 1617 176 1621 180
rect 1553 168 1557 172
rect 1537 160 1541 164
rect 1471 152 1475 156
rect 1455 144 1459 148
rect 1391 136 1395 140
rect 1375 128 1379 132
use shiftData  shiftData_1
timestamp 1749990304
transform 1 0 1312 0 1 218
box -4 166 1306 226
<< end >>
