magic
tech scmos
timestamp 1748092460
<< nwell >>
rect -1 -26 11 -15
<< polysilicon >>
rect 4 -20 6 -17
rect 4 -26 6 -24
<< pdiffusion >>
rect 3 -24 4 -20
rect 6 -24 7 -20
<< ptransistor >>
rect 4 -24 6 -20
<< polycontact >>
rect 3 -17 7 -13
<< pdcontact >>
rect -1 -24 3 -20
rect 7 -24 11 -20
<< end >>
