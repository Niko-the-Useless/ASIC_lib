magic
tech scmos
timestamp 1748092460
<< pwell >>
rect -132 -49 -118 -29
<< nwell >>
rect -132 -19 -107 -7
<< metal1 >>
rect -127 -11 -113 -7
rect -134 -37 -130 -11
rect -127 -19 -113 -15
rect -127 -33 -123 -19
rect -110 -41 -106 -11
rect -120 -45 -106 -41
use nmos  nmos_0
timestamp 1748092009
transform 0 -1 -145 -1 0 -32
box -3 -24 9 -11
use nmos  nmos_1
timestamp 1748092009
transform 0 1 -105 -1 0 -40
box -3 -24 9 -11
use pmos  pmos_0
timestamp 1748092460
transform 0 -1 -147 -1 0 -8
box -1 -26 11 -13
use pmos  pmos_1
timestamp 1748092460
transform 0 1 -93 -1 0 -8
box -1 -26 11 -13
<< labels >>
rlabel pwell -127 -49 -123 -45 1 Gnd
rlabel metal1 -127 -11 -113 -7 5 Vdd
rlabel metal1 -134 -37 -130 -11 3 A
rlabel metal1 -127 -33 -123 -15 1 NAND
rlabel metal1 -110 -45 -106 -11 7 B
<< end >>
