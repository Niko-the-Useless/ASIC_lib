magic
tech scmos
timestamp 1749993027
<< pwell >>
rect -19 -44 33 -32
<< nwell >>
rect -19 -22 33 -10
<< polysilicon >>
rect -14 -15 -12 -4
rect -6 -15 -4 -4
rect 2 -15 4 -4
rect 10 -15 12 -4
rect 24 -17 27 -15
rect 31 -17 33 -15
rect -14 -36 -12 -18
rect -6 -36 -4 -18
rect 2 -36 4 -18
rect 10 -36 12 -18
rect -14 -44 -12 -39
rect -6 -44 -4 -39
rect 2 -44 4 -39
rect 10 -44 12 -39
rect 24 -39 27 -37
rect 31 -39 33 -37
<< ndiffusion >>
rect -15 -39 -14 -36
rect -12 -39 -11 -36
rect -7 -39 -6 -36
rect -4 -39 -3 -36
rect 1 -39 2 -36
rect 4 -39 5 -36
rect 9 -39 10 -36
rect 12 -39 13 -36
rect 27 -37 31 -36
rect 27 -40 31 -39
<< pdiffusion >>
rect -15 -18 -14 -15
rect -12 -18 -11 -15
rect -7 -18 -6 -15
rect -4 -18 -3 -15
rect 1 -18 2 -15
rect 4 -18 5 -15
rect 9 -18 10 -15
rect 12 -18 13 -15
rect 27 -15 31 -14
rect 27 -18 31 -17
<< metal1 >>
rect -25 -10 31 -7
rect -25 -11 27 -10
rect -19 -14 -15 -11
rect -3 -14 1 -11
rect 13 -14 17 -11
rect -11 -25 -7 -18
rect 5 -25 9 -18
rect 20 -25 24 -18
rect -19 -29 24 -25
rect 13 -36 17 -29
rect 20 -36 24 -29
rect 27 -32 31 -22
rect -19 -43 -15 -40
rect -19 -44 27 -43
rect -19 -47 31 -44
<< ntransistor >>
rect -14 -39 -12 -36
rect -6 -39 -4 -36
rect 2 -39 4 -36
rect 10 -39 12 -36
rect 27 -39 31 -37
<< ptransistor >>
rect -14 -18 -12 -15
rect -6 -18 -4 -15
rect 2 -18 4 -15
rect 10 -18 12 -15
rect 27 -17 31 -15
<< polycontact >>
rect -15 -4 -11 0
rect -7 -4 -3 0
rect 1 -4 5 0
rect 9 -4 13 0
rect 20 -18 24 -14
rect 20 -40 24 -36
<< ndcontact >>
rect 27 -36 31 -32
rect -19 -40 -15 -36
rect -11 -40 -7 -36
rect -3 -40 1 -36
rect 5 -40 9 -36
rect 13 -40 17 -36
rect 27 -44 31 -40
<< pdcontact >>
rect -19 -18 -15 -14
rect -11 -18 -7 -14
rect -3 -18 1 -14
rect 5 -18 9 -14
rect 27 -14 31 -10
rect 13 -18 17 -14
rect 27 -22 31 -18
<< end >>
