magic
tech scmos
timestamp 1749982892
<< metal1 >>
rect 1297 436 1333 440
rect 1296 391 1332 395
rect 19 376 2625 380
rect 19 368 2598 372
rect 2602 368 2625 372
rect 19 360 2534 364
rect 2538 360 2625 364
rect 19 352 2518 356
rect 2522 352 2625 356
rect 19 344 2452 348
rect 2456 344 2625 348
rect 19 336 2436 340
rect 2440 336 2625 340
rect 19 328 2372 332
rect 2376 328 2625 332
rect 19 320 2356 324
rect 2360 320 2625 324
rect 19 312 2287 316
rect 2291 312 2625 316
rect 19 304 2271 308
rect 2275 304 2625 308
rect 19 296 2207 300
rect 2211 296 2625 300
rect 19 288 2191 292
rect 2195 288 2625 292
rect 19 280 2125 284
rect 2129 280 2625 284
rect 19 272 2109 276
rect 2113 272 2625 276
rect 19 264 2045 268
rect 2049 264 2625 268
rect 19 256 2029 260
rect 2033 256 2625 260
rect 19 248 1960 252
rect 1964 248 2625 252
rect 19 240 1944 244
rect 1948 240 2625 244
rect 19 232 1880 236
rect 1884 232 2625 236
rect 19 224 1864 228
rect 1868 224 2625 228
rect 19 216 1798 220
rect 1802 216 2625 220
rect 19 208 1782 212
rect 1786 208 2625 212
rect 19 200 1718 204
rect 1722 200 2625 204
rect 19 192 1702 196
rect 1706 192 2625 196
rect 19 184 1633 188
rect 1637 184 2625 188
rect 19 176 1617 180
rect 1621 176 2625 180
rect 19 168 1553 172
rect 1557 168 2625 172
rect 19 160 1537 164
rect 1541 160 2625 164
rect 19 152 1471 156
rect 1475 152 2625 156
rect 19 144 1455 148
rect 1459 144 2625 148
rect 19 136 1391 140
rect 1395 136 2625 140
rect 19 128 1375 132
rect 1379 128 2625 132
rect 19 120 1306 124
rect 1310 120 2625 124
rect 19 112 1290 116
rect 1294 112 2625 116
rect 19 104 1226 108
rect 1230 104 2625 108
rect 19 96 1210 100
rect 1214 96 2625 100
rect 19 88 1144 92
rect 1148 88 2625 92
rect 19 80 1128 84
rect 1132 80 2625 84
rect 19 72 1064 76
rect 1068 72 2625 76
rect 19 64 1048 68
rect 1052 64 2625 68
rect 19 56 979 60
rect 983 56 2625 60
rect 19 48 963 52
rect 967 48 2625 52
rect 19 40 899 44
rect 903 40 2625 44
rect 19 32 883 36
rect 887 32 2625 36
rect 19 24 817 28
rect 821 24 2625 28
rect 19 16 801 20
rect 805 16 2625 20
rect 19 8 737 12
rect 741 8 2625 12
rect 19 0 721 4
rect 725 0 2625 4
rect 19 -8 652 -4
rect 656 -8 2625 -4
rect 19 -16 636 -12
rect 640 -16 2625 -12
rect 19 -24 572 -20
rect 576 -24 2625 -20
rect 19 -32 556 -28
rect 560 -32 2625 -28
rect 19 -40 490 -36
rect 494 -40 2625 -36
rect 19 -48 474 -44
rect 478 -48 2625 -44
rect 19 -56 410 -52
rect 414 -56 2625 -52
rect 19 -64 394 -60
rect 398 -64 2625 -60
rect 19 -72 325 -68
rect 329 -72 2625 -68
rect 19 -80 309 -76
rect 313 -80 2625 -76
rect 19 -88 245 -84
rect 249 -88 2625 -84
rect 19 -96 229 -92
rect 233 -96 2625 -92
rect 19 -104 163 -100
rect 167 -104 2625 -100
rect 19 -112 147 -108
rect 151 -112 2625 -108
rect 19 -120 83 -116
rect 87 -120 2625 -116
rect 19 -128 67 -124
rect 71 -128 2625 -124
<< metal2 >>
rect 1266 440 1340 444
rect 67 -124 71 388
rect 83 -116 87 388
rect 147 -108 151 388
rect 163 -100 167 388
rect 229 -92 233 388
rect 245 -84 249 388
rect 309 -76 313 388
rect 325 -68 329 388
rect 394 -60 398 388
rect 410 -52 414 388
rect 474 -44 478 388
rect 490 -36 494 388
rect 556 -28 560 388
rect 572 -20 576 388
rect 636 -12 640 388
rect 652 -4 656 388
rect 721 4 725 388
rect 737 12 741 388
rect 801 20 805 388
rect 817 28 821 388
rect 883 36 887 388
rect 899 44 903 388
rect 963 52 967 388
rect 979 60 983 388
rect 1048 68 1052 388
rect 1064 76 1068 388
rect 1128 84 1132 388
rect 1144 92 1148 388
rect 1210 100 1214 388
rect 1226 108 1230 388
rect 1290 116 1294 419
rect 1306 124 1310 419
rect 1375 132 1379 388
rect 1391 140 1395 388
rect 1455 148 1459 388
rect 1471 156 1475 388
rect 1537 164 1541 388
rect 1553 172 1557 388
rect 1617 180 1621 388
rect 1633 188 1637 388
rect 1702 196 1706 388
rect 1718 204 1722 388
rect 1782 212 1786 388
rect 1798 220 1802 388
rect 1864 228 1868 388
rect 1880 236 1884 388
rect 1944 244 1948 388
rect 1960 252 1964 388
rect 2029 260 2033 388
rect 2045 268 2049 388
rect 2109 276 2113 399
rect 2125 284 2129 399
rect 2191 292 2195 419
rect 2207 300 2211 419
rect 2271 308 2275 392
rect 2287 316 2291 392
rect 2356 324 2360 392
rect 2372 332 2376 392
rect 2436 340 2440 392
rect 2452 348 2456 392
rect 2518 356 2522 392
rect 2534 364 2538 392
rect 2598 372 2602 392
rect 2614 376 2618 393
<< m2contact >>
rect 2598 368 2602 372
rect 2534 360 2538 364
rect 2518 352 2522 356
rect 2452 344 2456 348
rect 2436 336 2440 340
rect 2372 328 2376 332
rect 2356 320 2360 324
rect 2287 312 2291 316
rect 2271 304 2275 308
rect 2207 296 2211 300
rect 2191 288 2195 292
rect 2125 280 2129 284
rect 2109 272 2113 276
rect 2045 264 2049 268
rect 2029 256 2033 260
rect 1960 248 1964 252
rect 1944 240 1948 244
rect 1880 232 1884 236
rect 1864 224 1868 228
rect 1798 216 1802 220
rect 1782 208 1786 212
rect 1718 200 1722 204
rect 1702 192 1706 196
rect 1633 184 1637 188
rect 1617 176 1621 180
rect 1553 168 1557 172
rect 1537 160 1541 164
rect 1471 152 1475 156
rect 1455 144 1459 148
rect 1391 136 1395 140
rect 1375 128 1379 132
rect 1306 120 1310 124
rect 1290 112 1294 116
rect 1226 104 1230 108
rect 1210 96 1214 100
rect 1144 88 1148 92
rect 1128 80 1132 84
rect 1064 72 1068 76
rect 1048 64 1052 68
rect 979 56 983 60
rect 963 48 967 52
rect 899 40 903 44
rect 883 32 887 36
rect 817 24 821 28
rect 801 16 805 20
rect 737 8 741 12
rect 721 0 725 4
rect 652 -8 656 -4
rect 636 -16 640 -12
rect 572 -24 576 -20
rect 556 -32 560 -28
rect 490 -40 494 -36
rect 474 -48 478 -44
rect 410 -56 414 -52
rect 394 -64 398 -60
rect 325 -72 329 -68
rect 309 -80 313 -76
rect 245 -88 249 -84
rect 229 -96 233 -92
rect 163 -104 167 -100
rect 147 -112 151 -108
rect 83 -120 87 -116
rect 67 -128 71 -124
use shiftData  shiftData_0
timestamp 1749982892
transform 1 0 4 0 1 218
box -4 166 1306 235
use shiftData  shiftData_1
timestamp 1749982892
transform 1 0 1312 0 1 218
box -4 166 1306 235
<< end >>
