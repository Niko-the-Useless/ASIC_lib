magic
tech scmos
timestamp 1748362390
<< pwell >>
rect -20 -20 -9 -8
<< nwell >>
rect -20 2 -9 14
<< polysilicon >>
rect -18 7 -15 9
rect -11 7 -9 9
rect -18 -15 -15 -13
rect -11 -15 -9 -13
<< ndiffusion >>
rect -15 -13 -11 -12
rect -15 -16 -11 -15
<< pdiffusion >>
rect -15 9 -11 10
rect -15 6 -11 7
<< metal1 >>
rect -22 -12 -18 6
rect -15 -8 -11 2
<< ntransistor >>
rect -15 -15 -11 -13
<< ptransistor >>
rect -15 7 -11 9
<< polycontact >>
rect -22 6 -18 10
rect -22 -16 -18 -12
<< ndcontact >>
rect -15 -12 -11 -8
rect -15 -20 -11 -16
<< pdcontact >>
rect -15 10 -11 14
rect -15 2 -11 6
<< end >>
