magic
tech scmos
timestamp 1748090986
<< pwell >>
rect -8 -20 3 -8
<< nwell >>
rect -8 2 3 14
<< polysilicon >>
rect -6 7 -3 9
rect 1 7 3 9
rect -6 -15 -3 -13
rect 1 -15 3 -13
<< ndiffusion >>
rect -3 -13 1 -12
rect -3 -16 1 -15
<< pdiffusion >>
rect -3 9 1 10
rect -3 6 1 7
<< metal1 >>
rect -3 14 1 18
rect -10 -1 -6 6
rect -15 -5 -6 -1
rect -10 -12 -6 -5
rect -3 -1 1 2
rect -3 -5 6 -1
rect -3 -8 1 -5
rect -3 -24 1 -20
<< ntransistor >>
rect -3 -15 1 -13
<< ptransistor >>
rect -3 7 1 9
<< polycontact >>
rect -10 6 -6 10
rect -10 -16 -6 -12
<< ndcontact >>
rect -3 -12 1 -8
rect -3 -20 1 -16
<< pdcontact >>
rect -3 10 1 14
rect -3 2 1 6
<< labels >>
rlabel metal1 -15 -5 -6 -1 3 A
rlabel metal1 -3 -24 1 -20 1 Gnd
rlabel metal1 -3 14 1 18 5 Vdd
rlabel metal1 -3 -5 6 -1 7 NA
<< end >>
