magic
tech scmos
timestamp 1742802863
<< checkpaint >>
rect 16 -3 34 11
<< nwell >>
rect 17 -2 33 8
<< polysilicon >>
rect 24 6 26 7
rect 24 -3 26 0
<< pdiffusion >>
rect 17 5 24 6
rect 20 1 24 5
rect 17 0 24 1
rect 26 5 33 6
rect 26 1 30 5
rect 26 0 33 1
<< ptransistor >>
rect 24 0 26 6
<< polycontact >>
rect 23 7 27 11
<< pdcontact >>
rect 16 1 20 5
rect 30 1 34 5
<< labels >>
rlabel pdcontact 16 1 20 5 1 source
rlabel pdcontact 30 1 34 5 7 drain
rlabel polycontact 23 7 27 11 5 gate
<< end >>
