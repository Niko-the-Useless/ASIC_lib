magic
tech scmos
timestamp 1749990304
<< metal1 >>
rect 158 52 188 56
rect 158 7 187 11
<< metal2 >>
rect 27 56 31 60
rect 123 56 193 60
use shiftreg2  shiftreg2_0
timestamp 1749982892
transform 1 0 0 0 1 7
box 0 -7 167 53
use shiftreg2  shiftreg2_1
timestamp 1749982892
transform 1 0 162 0 1 7
box 0 -7 167 53
<< end >>
